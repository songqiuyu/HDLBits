module top_module (
    input clk,
    input areset,
    input x,
    output z
); 

    //Mealy
    // Implement using one-hot encoding. 



endmodule