//no input, one output 输出一个1
module top_module( output one);
	assign one = 1;
endmodule