//实现二维元胞自动机
            /**
            0   [0:15]
            1   [16:31]
            2   [32:47]
            3   [48:63]
            4   64
            5   80
            6   16*6
            7   16*7
            8
            9
            10
            11
            12
            13
            14
            15
            **/
module top_module(
    input clk,
    input load,
    input [255:0] data,
    output reg [255:0] q ); 
// Hint中提示边界检测
    integer i, j;
    integer t;
    always@(posedge clk)begin
        if(load)
            q <= data;
        else begin
        /**
                当前行列为 i, j
                上方，行-1，列不变  ((i-1+16)%16)*16 + j
                下方，行+1，列不变  ((i+1)%16)*16 + j
                左方，行不变，列-1  i*16 + (j-1+16)%16
                右方，行不变，列+1  i*16 + (j+1)%16
                左上方，行-1，列-1  ((i-1+16)%16)*16 + (j-1+16)%16
                右上方，行-1，列+1  ((i-1+16)%16)*16 + (j+1)%16
                左下方，行+1，列-1  ((i+1)%16)*16 + (j-1+16)%16
                右下方，行+1，列+1  ((i+1)%16)*16 + (j+1)%16

        **/

        // 要注意区分阻塞和非阻塞，t就不能用非阻塞！

            for(i=0;i<=15;i=i+1)begin
                for(j=0;j<=15;j=j+1)begin
                    //一定是=而不是<=
                    t = q[((i-1+16)%16)*16 + j] + q[((i+1)%16)*16 + j] + q[i*16 + (j-1+16)%16] + q[i*16 + (j+1)%16] + q[((i-1+16)%16)*16 + (j-1+16)%16] + q[((i-1+16)%16)*16 + (j+1)%16] + q[((i+1)%16)*16 + (j-1+16)%16] + q[((i+1)%16)*16 + (j+1)%16];
                    if(t < 2 || t >3)
                        q[i*16 + j] <= 0;
                    else if(t == 3)
                        q[i*16 + j] <= 1; 
                end
            end
        end
    

    end


endmodule