//Create a module that implements a NOT gate.
// ~表示取反 
module top_module( input in, output out );
	assign out = ~in;
endmodule