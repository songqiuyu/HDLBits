//the ripple carry adder
//���мӷ��������мӷ����ڶ�������Ҫ�ȵ�һ�������ٽ��м���
//carry-select adder�ǽ�λѡ��ӷ���

module top_module(

);

endmodule

module add16 ( 
    input[15:0] a, 
    input[15:0] b, 
    input cin, 
    output[15:0] sum, 
    output cout );



endmodule